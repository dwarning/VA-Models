transient test circuit for igbt model 

.model my_igbt igbt3

va Vaa 0 dc 300
LL Vaa 1 80u
RL 1 a 30
Yigbt3 igbt1 a g 0 my_igbt
vg gg 0 PULSE(0 20 20us 100ns 100ns 50us 100us)
Rg gg g 100

.tran 10n 100u
.print tran v(g) V(a)
.end
