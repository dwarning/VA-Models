EKV 3.02 dioden test

.include ../Modelcards/90nm_xyce.lib

vd  d 0 dc 0.0
vg  g 0 dc 0.0
vs  s 0 dc 0.0
vb  b 0 dc 0.0
Yekv3_rf m1 d g s b pmos90 W=5e-6 L=0.5e-6

.dc vb 3 -0.1 -0.01 temp -50 150 50
.print dc i(vd)

.end

