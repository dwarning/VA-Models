Sample netlist BSIM6: Id plot nmos

.include "../Modelcards/modelcard_va.nmos"

vd d 0 dc 50m
vg g 0 dc 0.0
vs s 0 dc 0.0
vb b 0 dc 0.0

Ybsim6_va m1 d g s b nmos W = 10e-6 L = 1e-6

.step vb 0.0 -0.5 -0.1
.dc vg 0.0 1.2 0.01
.print dc format=gnuplot v(g) i(vd)
*.dc vd 0.0 1.2 0.01 vg 0.4 1.0 0.3
*.print dc v(d) i(vd)

.end

