ECL DFF HICUM2.4 test case
*
V6 D 0 dc 0 PULSE(-.25 0 0 1P 1P .25N .50N)   
V5 D_BAR 0 dc 0 PULSE(0 -.25 0 1P 1P .25N .50N)   
V4 CLK 0 dc 0 PULSE(-0.9 -1.2 0 1P 1P .125N .25N)   
V3 CLK_BAR 0 dc 0 PULSE(-1.2 -0.9 0 1P 1P .125N .25N)   
VVCS NET2 0 DC -0.8 
R6 0 NET6  800 
R5 0 NET11  800 
R4 NET12 VEE  350 
VVEE VEE 0 DC -2.0 
R3 0 NET10  800 
R2 NET13 VEE  350 
R1 0 Q  800 
XQVLGNPN16 NET7 CLK_BAR NET4 VEE dt hicumL0V1p1_c_sbt
XQVLGNPN15 NET5 CLK NET3 VEE dt hicumL0V1p1_c_sbt
XQVLGNPN14 NET1dt Q NET7 VEE dt hicumL0V1p1_c_sbt
XQVLGNPN13 Q NET6 NET9 VEE dt hicumL0V1p1_c_sbt
XQVLGNPN12 NET6 NET11 NET5 VEE dt hicumL0V1p1_c_sbt
XQVLGNPN11 NET11 D_BAR NET8 VEE dt hicumL0V1p1_c_sbt
XQVLGNPN1dt NET4 NET2 NET13 VEE dt hicumL0V1p1_c_sbt
XQVLGNPN9 NET3 NET2 NET12 VEE dt hicumL0V1p1_c_sbt
XQVLGNPN8 NET8 CLK_BAR NET3 VEE dt hicumL0V1p1_c_sbt
XQVLGNPN7 NET9 CLK NET4 VEE dt hicumL0V1p1_c_sbt
XQVLGNPN6 Q NET1dt NET7 VEE dt hicumL0V1p1_c_sbt
XQVLGNPN5 NET1dt NET11 NET9 VEE dt hicumL0V1p1_c_sbt
XQVLGNPN4 NET11 NET6 NET5 VEE dt hicumL0V1p1_c_sbt
XQVLGNPN3 NET6 D NET8 VEE dt hicumL0V1p1_c_sbt

Rdt dt 0 1G
*
.include ../Modelcards/model-card-hicumL0V1p11_mod_X.lib
.TRAN 0.25p 5n
.print tran format=gnuplot V(D) V(CLK) V(Q)

.END
