** One-Bit Comparator (Tran): Benchmarking Implementation of BSIM4.8.0 

Ybsim4va M1 Anot A Vdd Vdd P1  W=3.6u L=0.2u
Ybsim4va M2 Anot A 0 0 N1 W=1.8u L=0.2u
Ybsim4va M3 Bnot B Vdd Vdd  P1 W=3.6u L=0.2u
Ybsim4va M4 Bnot B 0 0 N1 W=1.8u L=0.2u
Ybsim4va M5 AorBnot 0 Vdd Vdd P1 W=1.8u L=3.6u
Ybsim4va M6 AorBnot B 1 0 N1 W=1.8u L=0.2u
Ybsim4va M7 1 Anot 0 0 N1 W=1.8u L=0.2u
Ybsim4va M8 Lnot 0 Vdd Vdd P1 W=1.8u L=3.6u
Ybsim4va M9 Lnot Bnot 2 0 N1 W=1.8u L=0.2u
Ybsim4va M10 2 A 0 0 N1 W=1.8u L=0.2u
Ybsim4va M11 Qnot 0 Vdd Vdd P1 W=3.6u L=3.6u
Ybsim4va M12 Qnot AorBnot 3 0 N1 W=1.8u L=0.2u
Ybsim4va M13 3 Lnot 0 0 N1 W=1.8u L=0.2u
Ybsim4va MQLO 8 Qnot Vdd Vdd  P1 W=3.6u L=0.2u
Ybsim4va MQL1 8 Qnot 0 0 N1 W=1.8u L=0.2u
Ybsim4va MLTO 9 Lnot Vdd Vdd P1 W=3.6u L=0.2u
Ybsim4va MLT1 9 Lnot 0 0 N1 W=1.8u L=0.2u
CQ Qnot 0 30f
CL Lnot 0 10f

Vdd Vdd 0 1.8
Va A 0  pulse 0 1.8 10ns .1ns .1ns 15ns 30ns
Vb B 0 0

.include "../Modelcards/modelcard.nmos"
.include "../Modelcards/modelcard.pmos"

.tran 1ns 60ns
.print tran v(a) v(b) v(9) v(8) 

.end
