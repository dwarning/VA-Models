Test of EKV3 noise

.include "../Modelcards/ekv3_150nm.mod"
Yekv3_rf M1 D G 0 0 NMOS150 W=150e-9 L=150e-9  NF=1

Vg G Ga DC .7v AC 1
Vgprobe 0 Ga 0
Vd 1 Da DC 1v
Ldrain 1 D 1
Cdrain D 0 1
*Rdrain 2 0 1
Vdprobe 0 Da 0

.options device temp=25
.noise V(D) vg dec 11 1k 100g 1
.print noise inoise onoise

* Verify that case does not matter in the device names or noise type names
* for the DNO and DNI operators.
*.print noise {sqrt(abs(inoise))} {pow(abs(onoise),1/3)}
*+ {pow(abs(DNO(M1,flicker_b_gnd)),1/3)}
*+ {pow(abs(DNO(M1,flicker_di_si_flicker_noise_in_channel_internal_nodes_#2)),1/3)}
*+ {pow(abs(DNO(M1,flicker_g_gnd_gate_flicker_noise)),1/3)}
*+ {pow(abs(DNO(M1,white_d_di)),1/3)}
*+ {pow(abs(DNO(M1,white_di_si)),1/3)}
*+ {pow(abs(DNO(M1,white_di_si_thermal_noise_in_channel_internal_nodes_#2)),1/3)}
*+ {pow(abs(DNO(M1,white_g_gnd_gate_shot_noise)),1/3)}
*+ {pow(abs(DNO(M1,white_noi_gnd)),1/3)}
*+ {pow(abs(DNO(M1,white_s_si)),1/3)}
*+ {pow(abs(DNO(m1)),1/3)}
*+ {pow(abs(DNI(M1,flicker_b_gnd)),1/3)}
*+ {pow(abs(DNI(M1,flicker_di_si_flicker_noise_in_channel_internal_nodes_#2)),1/3)}
*+ {pow(abs(DNI(M1,flicker_g_gnd_gate_flicker_noise)),1/3)}
**+ {pow(abs(DNI(M1,white_d_di)),1/3)}
*+ {pow(abs(DNI(M1,white_di_si)),1/3)}
*+ {pow(abs(DNI(M1,white_di_si_thermal_noise_in_channel_internal_nodes_#2)),1/3)}
*+ {pow(abs(DNI(M1,white_g_gnd_gate_shot_noise)),1/3)}
*+ {pow(abs(DNI(M1,white_noi_gnd)),1/3)}
**+ {pow(abs(DNI(M1,white_s_si)),1/3)}
*+ {pow(abs(DNI(m1)),1/3)}

.end
