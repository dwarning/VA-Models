** One-Shot Trigger (Tran): by Weidong Liu 5/16/2000.

yekv3_rf md1 4 in Vdd Vdd pmos90 W=0.36u L=0.12u ad=4e-12 as=4e-12
yekv3_rf md2 4 in 0 0 nmos90 W=0.18u L=0.12u ad=2e-12 as=2e-12
c4 4 0 30f
yekv3_rf md3 A 4 Vdd Vdd pmos90 W=0.36u L=0.12u ad=4e-12 as=4e-12
yekv3_rf md4 A 4 0 0 nmos90 W=0.18u L=0.12u ad=2e-12 as=2e-12
ca A 0 30f

yekv3_rf m1 Anot A Vdd Vdd pmos90 W=0.36u L=0.12u ad=4e-12 as=4e-12
yekv3_rf m2 Anot A 0 0 nmos90 W=0.18u L=0.12u ad=2e-12 as=2e-12

yekv3_rf m3 Bnot in Vdd Vdd pmos90 W=0.36u L=0.12u ad=4e-12 as=4e-12
yekv3_rf m4 Bnot in 0 0 nmos90 W=0.18u L=0.12u ad=2e-12 as=2e-12

yekv3_rf m5 AorBnot 0 Vdd Vdd pmos90 W=0.18u L=0.36u ad=2e-12 as=2e-12
yekv3_rf m6 AorBnot in 1 0 nmos90 W=0.18u L=0.12u ad=2e-12 as=2e-12
yekv3_rf m7 1 Anot 0 0 nmos90 W=0.18u L=0.12u ad=2e-12 as=2e-12

yekv3_rf m8 Lnot 0 Vdd Vdd pmos90 W=0.18u L=0.36u ad=4e-12 as=4e-12
yekv3_rf m9 Lnot Bnot 2 0 nmos90 W=0.18u L=0.12u ad=2e-12 as=2e-12
yekv3_rf m10 2 A 0 0 nmos90 W=0.18u L=0.12u ad=2e-12 as=2e-12

yekv3_rf m11 out 0 Vdd Vdd pmos90 W=0.36u L=0.36u ad=4e-12 as=4e-12
yekv3_rf m12 out AorBnot 3 0 nmos90 W=0.18u L=0.12u ad=2e-12 as=2e-12
yekv3_rf m13 3 Lnot 0 0 nmos90 W=0.18u L=0.12u ad=2e-12 as=2e-12

Vcc Vdd 0 1.8
vin in 0 pulse(0 1.8 1ns .1ns .1ns .8ns 5ns)

.tran .1ns 10ns
.include ../Modelcards/90nm_xyce.lib

.print tran v(in) v(out)

.end