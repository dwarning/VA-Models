** One-Bit Comparator (Tran): by Weidong Liu 5/16/2000.

yekv26_va m1 Anot A Vdd Vdd  pch W=3.6u L=1.2u
yekv26_va m2 Anot A 0 0 nch W=1.8u L=1.2u
yekv26_va m3 Bnot B Vdd Vdd  pch W=3.6u L=1.2u
yekv26_va m4 Bnot B 0 0 nch W=1.8u L=1.2u
yekv26_va m5 AorBnot 0 Vdd Vdd pch W=1.8u L=3.6u
yekv26_va m6 AorBnot B 1 0 nch W=1.8u L=1.2u
yekv26_va m7 1 Anot 0 0 nch W=1.8u L=1.2u
yekv26_va m8 Lnot 0 Vdd Vdd pch W=1.8u L=3.6u
yekv26_va m9 Lnot Bnot 2 0 nch W=1.8u L=1.2u
yekv26_va m10 2 A 0 0 nch W=1.8u L=1.2u
yekv26_va m11 Qnot 0 Vdd Vdd pch W=3.6u L=3.6u
yekv26_va m12 Qnot AorBnot 3 0 nch W=1.8u L=1.2u
yekv26_va m13 3 Lnot 0 0 nch W=1.8u L=1.2u
yekv26_va mQLO 8 Qnot Vdd Vdd  pch W=3.6u L=1.2u
yekv26_va mQL1 8 Qnot 0 0 nch W=1.8u L=1.2u
yekv26_va mLTO 9 Lnot Vdd Vdd pch W=3.6u L=1.2u
yekv26_va mLT1 9 Lnot 0 0 nch W=1.8u L=1.2u
CQ Qnot 0 30f
CL Lnot 0 10f

Vdd Vdd 0 1.8
Va A 0  pulse 0 1.8 10ns .1ns .1ns 15ns 30ns
Vb B 0 0

.tran .1ns 60ns
.include ../Modelcards/ekv26_0u5.par

.print tran v(A) v(B) v(9) v(8)
.endc

.end