* Sample netlist: Id-Vd plot *

.include ../Modelcards/model.l

vd d 0 dc 1.3
vg g 0 dc 0
vs s 0 dc 0
vb b 0 dc 0

Ybsimbulk m1 d g s b nmos W=10e-6 L=10e-6

.step vg 0.4 1 0.3
.dc vd 0.0 1.3 0.01
.print dc format=gnuplot v(d) i(vd)
*.probe dc ids=par'-i(vd)'
*.probe dc gds=deriv(ids)
*.print dc par'ids' par'gds'

.end
