MEXTRAM Gummel Test Ic,b,s=f(Vc,Ib)


VB B 0 0.5
VC C 0 1.0
VS S 0 0.0

*.model BJTRF1 bjt504_va
*Ybjt504_va q1 C B 0 S BJTRF1

.model BJTRF1 bjt504t_va
Ybjt504t_va q1 C B 0 S dt BJTRF1

*.model BJTRF1 bjt505_va
*Ybjt505_va q1 C B 0 S BJTRF1

*.model BJTRF1 bjt505t_va
*Ybjt505t_va q1 C B 0 S dt BJTRF1

*RT dt 0 100

*.op
.dc vb 0.2 1.4 0.01
.print dc v(B) i(vc) i(vb) i(vs)

.end
