dc test circuit for igbt model 

.model my_igbt igbt3

vg g 0 dc 10
vc a 0 dc 5
Yigbt3 igbt1 a g 0 my_igbt

.step vg 12.0 20.0 2.0
.dc vc 0.0 20.0 0.1
.print dc format=gnuplot v(g) v(a) i(vc)
.end