HICUM0 Gummel Test Ic=f(Vc,Vb)

VB B 0 0.5
VC C 0 1.0
VS S 0 0.0
XQ1 C B 0 S DT hicumL0V1p1_c_sbt
Rdt dt 0 10k

.dc vb 0.2 1.4 0.01
.print dc format=gnuplot v(b) i(vc) i(vb) i(vs)

.include ../Modelcards/model-card-hicumL0V1p11_mod_X.lib

.end
