Sample netlist for BSIM6
*Inverter Transient

.include "../Modelcards/modelcard.nmos"
.include "../Modelcards/modelcard.pmos"

* --- Voltage Sources ---
vdd   supply  0 dc 1.0
vin  vi  0 dc 0.5 sin (0.5 0.5 1MEG)

* --- Inverter Subcircuit ---
.subckt inverter vin vout vdd gnd
Ybsim6_va m1 vout vin vdd vdd pmos W = 20e-6 L = 1e-6
Ybsim6_va m2 vout vin gnd gnd nmos W = 10e-6 L = 1e-6
.ends

* --- Inverter ---
Xinv1  vi 1 supply 0 inverter
Xinv2  1 2 supply 0 inverter
Xinv3  2 3 supply 0 inverter
Xinv4  3 4 supply 0 inverter
Xinv5  4 vo supply 0 inverter

* --- Transient Analysis ---
.tran 10n 5u
.print tran v(vi) v(vo)

.end
