HICUM2v2.40 Gummel Test invers Ie,b,s=f(Ve,Ib) Vec=1V

VB B 0 1.2
VE E 0 1.0
VS S 0 0.0

YhicumL2_va q1 0 B E S dt hicumL2va
Rth dt 0 1.0

.dc vb 0.4 1.2 0.01
.print dc format=gnuplot v(b) i(ve) i(vb) i(vs)

.include ../Modelcards/examples_va.lib

.end
