Id-Vd Characteristics for L_UTSOI PMOS 

.model pmos1 l_utsoi_va type=-1

* --- Voltage Sources ---
vd drain 0 dc -0.05
vg gate 0 dc 1
vs source 0 dc 0
ve substrate 0 0

* --- Transistor ---
Yl_utsoi_va m1 drain gate source substrate tnode pmos1 W=1e-6 L=1e-7
*Yl_utsoi_va m1 drain gate source substrate pmos1 W=1e-6 L=1e-7
*Yl_utsoi_va m1 drain gate source substrate pmos1 W=1e-6 L=1e-7
*Yl_utsoi_va m1 drain gate source substrate 0 0 t pmos1 W=1e-6 L=1e-7

* --- DC Analysis ---
.dc vg -1.2 0.0 0.01
.print dc v(gate) i(vd)
*.dc vd -1.2 0 0.01 vg -1.2 -0.5 0.1
*.print dc i(vd)
*.print dc v(t)

.end
