Sample netlist for BSIMBULK
*Drain current symmetry for nmos

.include ../Modelcards/model.l

* --- Voltage Sources ---
vdrain drain 0 dc 0.0
esource source 0 drain 0 -1
vgate gate  0 dc 1.0
vbulk bulk 0 dc 0.0


* --- Transistor ---
Ybsimbulk m1 drain gate source bulk nmos W = 10e-6 L = 10e-6

* --- DC Analysis ---
.dc vdrain -0.1 0.1 0.001 vgate 0.0 1.0 0.2
.print dc i(vdrain)
*let gx=deriv(-i(vdrain))
*let gx2=deriv(gx)
*let gx3=deriv(gx2)
*plot gx
*plot gx2
*plot gx3

.end
