Bip model in subckt Gummel Test Ic=f(Vc,Vb)

VB B 0 0.5
VC C 0 1.0
VS S 0 0.0
X1 C B 0 S T bip_default

.dc vb 0.35 1.2 0.01
.print dc format=gnuplot i(vc) i(vb) i(vs)

********************************************************************************
* Complete test transistor: default
********************************************************************************
.subckt bip_default c b e s dt
YhicumL0va q1 c b e s dt hic0_full
.model hic0_full hicumL0va
.ends bip_default
********************************************************************************

.end
