Sample netlist for BSIMSOI
*17-stage ring oscillator

.include "../Modelcards/modelcard.nmos"
.include "../Modelcards/modelcard.pmos"

* --- Voltage Sources ---
vdd supply  0 dc 1.0

* --- Inverter Subcircuit ---
.subckt inverter vin vout vdd gnd
Ybsimsoi_va m1 vout vin vdd vdd pmos1 W = 20e-6 L = 1e-6
Ybsimsoi_va m2 vout vin gnd gnd nmos1 W = 10e-6 L = 1e-6
.ends

* --- 17 Stage Ring oscillator ---
Xinv1   1  2 supply 0 inverter
Xinv2   2  3 supply 0 inverter
Xinv3   3  4 supply 0 inverter
Xinv4   4  5 supply 0 inverter
Xinv5   5  6 supply 0 inverter
Xinv6   6  7 supply 0 inverter
Xinv7   7  8 supply 0 inverter
Xinv8   8  9 supply 0 inverter
Xinv9   9 10 supply 0 inverter
Xinv10 10 11 supply 0 inverter
Xinv11 11 12 supply 0 inverter
Xinv12 12 13 supply 0 inverter
Xinv13 13 14 supply 0 inverter
Xinv14 14 15 supply 0 inverter
Xinv15 15 16 supply 0 inverter
Xinv16 16 17 supply 0 inverter
Xinv17 17  1 supply 0 inverter

* --- Initial Condition ---
.ic  v(1)=1

.tran 1n 1u
.print tran v(1) v(17)

.end


