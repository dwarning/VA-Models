ECL DFF MEXTRAM test case
*
V6 D     GND PULSE(-.25 0 0 1P 1P .25N .50N)
V5 D_BAR GND PULSE(0 -.25 0 1P 1P .25N .50N)
V4 CLK     GND PULSE(-0.9 -1.2 0 1P 1P .125N .25N)
V3 CLK_BAR GND PULSE(-1.2 -0.9 0 1P 1P .125N .25N)
VVCS NET2 GND DC -0.8
R6 GND NET6  800
R5 GND NET11  800
R4 NET12 VEE  350
VEE VEE GND DC -2.0
R3 GND NET10  800
R2 NET13 VEE  350
R1 GND Q  800
NQVLGNPN16 NET7 CLK_BAR NET4 VEE BJTRF1
NQVLGNPN15 NET5 CLK NET3 VEE BJTRF1
NQVLGNPN14 NET10 Q NET7 VEE BJTRF1
NQVLGNPN13 Q NET6 NET9 VEE BJTRF1
NQVLGNPN12 NET6 NET11 NET5 VEE BJTRF1
NQVLGNPN11 NET11 D_BAR NET8 VEE BJTRF1
NQVLGNPN10 NET4 NET2 NET13 VEE BJTRF1
NQVLGNPN9 NET3 NET2 NET12 VEE BJTRF1
NQVLGNPN8 NET8 CLK_BAR NET3 VEE BJTRF1
NQVLGNPN7 NET9 CLK NET4 VEE BJTRF1
NQVLGNPN6 Q NET10 NET7 VEE BJTRF1
NQVLGNPN5 NET10 NET11 NET9 VEE BJTRF1
NQVLGNPN4 NET11 NET6 NET5 VEE BJTRF1
NQVLGNPN3 NET6 D NET8 VEE BJTRF1

*.model BJTRF1 bjt504va
.model BJTRF1 bjt504tva
*.model BJTRF1 bjt505_va
*.model BJTRF1 bjt505t_va

.SAVE V(D) V(CLK) V(Q)
.control
*pre_osdi ../osdilibs/bjt504.osdi
pre_osdi ../osdilibs/bjt504t.osdi
*pre_osdi ../osdilibs/bjt505.osdi
*pre_osdi ../osdilibs/bjt505t.osdi
*op
TRAN 0.25p 10n
plot V(D) V(CLK) V(Q)
.endc
.END
