HICUM0 Output Test Ic=f(Vc,Ib)

IB 0 B 200n
VC C 0 2.0
VS S 0 0.0
*IB B 0 200n
*VC 0 C 2.0
*VS S 0 0.0
X1 C B 0 S DT hicumL0V1p1_c_sbt

Rdt dt 0 1G

.step ib 10u 100u 10u
.dc vc 0.0 3.0 0.05
.print dc format=gnuplot v(c) i(vc) v(dt)

.include ../Modelcards/model-card-hicumL0V1p11_mod_X.lib 

.end
