test hys.va in DC, TRAN and Homotopy

.model H1 hys

V1 1 0 1 sin(0 0.7 1k)
NYhys 0 1 ns H1

.control
pre_osdi hys.osdi
* DC analysis
dc V1 -1 1 0.01
*.print dc V(1) I(V1) N(Yhys!H1_ns);N(Yhys!H1_ns) internal node ns of instance Yhys
plot I(V1) vs V(1) retraceplot 
*plot I(V1) vs V(ns) retraceplot 
* transient simulation
tran 1u 2m
plot I(V1) vs V(1) retraceplot 
*plot I(V1) vs V(ns) retraceplot 
.endc

.end
