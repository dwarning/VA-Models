** MOSFET Gain Stage (AC): Benchmarking Implementation of BSIM4.8.0 

Ybsim4va m1 d g 0 0 n1 L=0.09u W=4u
Rsource 1 g 100k
Rload d vdd 1k

Vdd vdd 0 1.8 
Vin 1 0 dc 0.8 ac 1

.ac dec 10 100 1000Meg 
.print ac vdb(d)

.include "../Modelcards/modelcard.nmos"

.end
