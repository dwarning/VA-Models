VBIC Gummel Test Ic=f(Vc,Ib)

.model my_vbic vbic13_4t_va

ib 0 b 1u
vc c 0 1.0
vs s 0 0.0
yvbic13_4t_va vbic1 c b 0 s my_vbic

.step ib 10u 100u 10u
.dc vc 0.0 5.0 0.01
.print dc format=gnuplot v(c) i(vc) i(vs)

.end
