Sample netlist BSIM6: Id plot pmos

.include "../Modelcards/modelcard_va.pmos"

vd d 0 dc -50m
vg g 0 dc 0.0
vs s 0 dc 0.0
vb b 0 dc 0.0

Ybsim6_va m1 d g s b pmos W = 20e-6 L = 1e-6

.step vb 0.0 0.5 0.1
.dc vg -1.2 0.0 0.01
.print dc format=gnuplot v(g) i(vd)
*.dc vd -1.2 0.0 0.01 vg -1.0 -0.4 0.2
*.print dc v(d) i(vd)

.end

