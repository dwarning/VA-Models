** One-Shot Trigger (Tran): Benchmarking Implementation of BSIM4.8.0 

Ybsim4va Md1 4 in Vdd Vdd  P1 W=3.6u L=0.2u
Ybsim4va Md2 4 in 0 0 N1 W=1.8u L=0.2u
c4 4 0 100f
Ybsim4va Md3 A 4 Vdd Vdd  P1 W=3.6u L=0.2u 
Ybsim4va Md4 A 4 0 0 N1 W=1.8u L=0.2u
ca a 0 100f

Ybsim4va M1 Anot A Vdd Vdd  P1 W=3.6u L=0.2u
Ybsim4va M2 Anot A 0 0 N1 W=1.8u L=0.2u

Ybsim4va M3 Bnot in Vdd Vdd  P1 W=3.6u L=0.2u
Ybsim4va M4 Bnot in 0 0 N1 W=1.8u L=0.2u

Ybsim4va M5 AorBnot 0 Vdd Vdd P1 W=1.8u L=3.6u
Ybsim4va M6 AorBnot in 1 0 N1 W=1.8u L=0.2u
Ybsim4va M7 1 Anot 0 0 N1 W=1.8u L=0.2u

Ybsim4va M8 Lnot 0 Vdd Vdd P1 W=1.8u L=3.6u
Ybsim4va M9 Lnot Bnot 2 0 N1 W=1.8u L=0.2u
Ybsim4va M10 2 A 0 0 N1 W=1.8u L=0.2u

Ybsim4va M11 out 0 Vdd Vdd P1 W=3.6u L=3.6u
Ybsim4va M12 out AorBnot 3 0 N1 W=1.8u L=0.2u
Ybsim4va M13 3 Lnot 0 0 N1 W=1.8u L=0.2u

Vcc vdd 0 1.8
vin in 0 pulse 0 1.8 1ns .1ns .1ns .8ns 5ns

.include "../Modelcards/modelcard.nmos"
.include "../Modelcards/modelcard.pmos"

.tran 1ns 10ns
.print tran v(in) v(out)

.end
