BSIMCMG Test

VD d 0 -0.05
VG g 0 -1
VS s 0 0
VB e 0 0

.include ../Modelcards/modelcard.pmos

Ybsimcmg_va m1 d g s e pmos L=0.2u NF=20

.step VG -0.5 -1.0 -0.1
.dc Vd 0 -1.0 -0.01
.print dc format=gnuplot v(d) i(VD)

.end
