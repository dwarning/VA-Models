r3_cmc

v1 1 0 10
Yr3_cmc r1 1 0 0 dt poly_87OhmPerSquare w=1.05u l=42u

* Poly resistor, r2_cmc model
.include ../Modelcards/poly_87OhmPerSquare.par

.step temp -40 160 40
.dc v1 -9.9 9.9 0.2
.print dc format=gnuplot v(1) '-v(1)/i(v1)'

.end
