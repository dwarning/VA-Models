* Sample netlist: Id-Vg plot *

.include ../Modelcards/model.l

vd d 0 dc -0.05
vg g 0 dc 0
vs s 0 dc 0
vb b 0 dc 0

Ybsimbulk m1 d g s b pmos W=10e-6 L=10e-6

.step vb 0 0.3 0.1
.dc vg -1.3 0.0 0.01
.print dc format=gnuplot v(g) i(vd)
*.probe dc ids=par'i(vd)'
*.probe dc gm=deriv(ids)
*.probe dc gm2=deriv(gm)
*.print dc par'ids' par'gm' par'gm2'

.end
