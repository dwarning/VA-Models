HICUM2v2.40 Output Test Ic=f(Vc,Ib)

IB 0 B 1u
VC C 0 1.8
VS S 0 0.0

YhicumL2_va q1 C B 0 S tj hicumL2va
rth tj 0 1g

.step ib 10u 100u 10u
.dc vc 0.0 1.8 0.01
.print dc format=gnuplot v(c) i(vc)
*.altermod @hicumL2va[flsh]=1
*.dc vc 0.0 1.8 0.01 ib 1u 10u 1u
*.plot -i(vc)
*.plot v(tj)

.include ../Modelcards/examples_va.lib

.end
