VBIC Gummel Test Ic=f(Vc,Vb)

.model my_vbic vbic13_4t_va

vb b 0 0.5
vc c 0 1.0
vs s 0 0.0
yvbic13_4t_va vbic1 c b 0 s my_vbic

.dc vb 0.2 1.2 0.01
.print dc v(b) i(vc) i(vb) i(vs)

.end
