Sample netlist for BSIMSOI

.include "../Modelcards/modelcard.nmos"

* --- Voltage Sources ---
vd d  0 dc 50m
vg g  0 dc 0.0
vs s  0 dc 0.0
vb b  0 dc 0.0

* --- Transistor ---
Ybsimsoi_va m1 d g s b nmos1 W = 10e-6 L = 1e-6

* --- DC Analysis ---
.step vb -0.5 0 0.1
.dc vg 0.0 1.2 0.01
.print dc format=gnuplot v(g) i(vd)
*.dc vd 0.0 1.2 0.01 vg 0.4 1.0 0.1
*.plot -i(vd)

.end

